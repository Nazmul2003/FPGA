----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Nazmul Haque
-- 
-- Create Date:    21:11:32 08/31/2023 
-- Design Name: 
-- Module Name:    primeBCD - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity primeBCD is
    Port ( A : in  STD_LOGIC_VECTOR (3 downto 0);
           f : out  STD_LOGIC);
end primeBCD;

architecture Behavioral of primeBCD is

begin

f <= (not A(3)) and ((A(2) and A(0)) or ((not A(2)) and A(1)));

end Behavioral;

